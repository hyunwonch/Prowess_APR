../../../../sim/DMA/dma_engine.sv