../../../../sim/PE_top/PE_array.sv