../../../../sim/Switch/switch.sv