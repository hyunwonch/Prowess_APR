../../../../sim/PE_top/PE_top.sv