`ifndef __PE_SVH__
`define __PE_SVH__

// word and register sizes
// typedef logic [31:0] ADDR;
// typedef logic [31:0] DATA;
// typedef logic [4:0] REG_IDX;
// typedef logic [63:0] INST;

// typedef struct packed {
//     logic [2:0] id,
//     INST inst2,
//     logic valid
// } CONTROL










`endif // __PE_SVH__