../../../../sim/DMA/dma.sv